module zk_stmt_arith(out, in);

output out;
input in;

assign out = in;

endmodule
